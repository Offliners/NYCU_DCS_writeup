module HE(
	// Input signals
	clk,
	rst_n,
	in_valid,
	in_image,
  // Output signals
	out_valid,
	out_image
);
//---------------------------------------------------------------------
//   INPUT AND OUTPUT DECLARATION                         
//---------------------------------------------------------------------
input				clk,rst_n,in_valid;
input [7:0]			in_image;
output logic 		out_valid;
output logic [7:0]	out_image;

//---------------------------------------------------------------------
// PARAMETER DECLARATION
//---------------------------------------------------------------------


//---------------------------------------------------------------------
//   LOGIC DECLARATION                             
//---------------------------------------------------------------------


//---------------------------------------------------------------------
//   Finite-State Mechine                                          
//---------------------------------------------------------------------


endmodule